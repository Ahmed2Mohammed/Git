module aa();

endmodule
